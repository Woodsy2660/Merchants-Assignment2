

module log10_lut (
    input [3:0] index,
    output reg [15:0] log10_value
);

always @(*) begin
    case (index)
        4'd0: log10_value = 16'd0;
        4'd1: log10_value = 16'd147;
        4'd2: log10_value = 16'd295;
        4'd3: log10_value = 16'd442;
        4'd4: log10_value = 16'd590;
        4'd5: log10_value = 16'd738;
        4'd6: log10_value = 16'd885;
        4'd7: log10_value = 16'd1033;
        4'd8: log10_value = 16'd1181;
        4'd9: log10_value = 16'd1328;
        4'd10: log10_value = 16'd1476;
        4'd11: log10_value = 16'd1624;
        4'd12: log10_value = 16'd1771;
        4'd13: log10_value = 16'd1919;
        4'd14: log10_value = 16'd2067;
        4'd15: log10_value = 16'd2214;
        default: log10_value = 16'd0;
    endcase
end

endmodule


