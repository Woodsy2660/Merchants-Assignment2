// vga.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module vga (
		input  wire       clk_clk,                     //           clk.clk
		input  wire [2:0] filter_select_filter_select, // filter_select.filter_select
		input  wire [7:0] intensity_intensity,         //     intensity.intensity
		input  wire [2:0] kernel_select_kernel_select, // kernel_select.kernel_select
		input  wire       reset_reset_n,               //         reset.reset_n
		output wire       vga_CLK,                     //           vga.CLK
		output wire       vga_HS,                      //              .HS
		output wire       vga_VS,                      //              .VS
		output wire       vga_BLANK,                   //              .BLANK
		output wire       vga_SYNC,                    //              .SYNC
		output wire [7:0] vga_R,                       //              .R
		output wire [7:0] vga_G,                       //              .G
		output wire [7:0] vga_B                        //              .B
	);

	wire         vga_face_0_avalon_streaming_source_valid;                           // vga_face_0:valid -> convolution_filter_wrapper_0:valid_in
	wire  [29:0] vga_face_0_avalon_streaming_source_data;                            // vga_face_0:data -> convolution_filter_wrapper_0:data_in
	wire         vga_face_0_avalon_streaming_source_ready;                           // convolution_filter_wrapper_0:ready_out -> vga_face_0:ready
	wire         vga_face_0_avalon_streaming_source_startofpacket;                   // vga_face_0:startofpacket -> convolution_filter_wrapper_0:startofpacket_in
	wire         vga_face_0_avalon_streaming_source_endofpacket;                     // vga_face_0:endofpacket -> convolution_filter_wrapper_0:endofpacket_in
	wire         convolution_filter_wrapper_0_avalon_streaming_source_valid;         // convolution_filter_wrapper_0:valid_out -> pixel_value_filter_0:valid_in
	wire  [29:0] convolution_filter_wrapper_0_avalon_streaming_source_data;          // convolution_filter_wrapper_0:data_out -> pixel_value_filter_0:data_in
	wire         convolution_filter_wrapper_0_avalon_streaming_source_ready;         // pixel_value_filter_0:ready_in -> convolution_filter_wrapper_0:ready_in
	wire         convolution_filter_wrapper_0_avalon_streaming_source_startofpacket; // convolution_filter_wrapper_0:startofpacket_out -> pixel_value_filter_0:startofpacket_in
	wire         convolution_filter_wrapper_0_avalon_streaming_source_endofpacket;   // convolution_filter_wrapper_0:endofpacket_out -> pixel_value_filter_0:endofpacket_in
	wire         pixel_value_filter_0_avalon_streaming_source_valid;                 // pixel_value_filter_0:valid_out -> video_vga_controller_0:valid
	wire  [29:0] pixel_value_filter_0_avalon_streaming_source_data;                  // pixel_value_filter_0:data_out -> video_vga_controller_0:data
	wire         pixel_value_filter_0_avalon_streaming_source_ready;                 // video_vga_controller_0:ready -> pixel_value_filter_0:ready_out
	wire         pixel_value_filter_0_avalon_streaming_source_startofpacket;         // pixel_value_filter_0:startofpacket_out -> video_vga_controller_0:startofpacket
	wire         pixel_value_filter_0_avalon_streaming_source_endofpacket;           // pixel_value_filter_0:endofpacket_out -> video_vga_controller_0:endofpacket
	wire         video_pll_0_vga_clk_clk;                                            // video_pll_0:vga_clk_clk -> [convolution_filter_wrapper_0:clk, pixel_value_filter_0:clk, rst_controller:clk, vga_face_0:clk, video_vga_controller_0:clk]
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [convolution_filter_wrapper_0:reset, pixel_value_filter_0:reset, vga_face_0:reset, video_vga_controller_0:reset]
	wire         video_pll_0_reset_source_reset;                                     // video_pll_0:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> video_pll_0:ref_reset_reset

	convolution_filter_wrapper #(
		.WIDTH  (640),
		.HEIGHT (480)
	) convolution_filter_wrapper_0 (
		.clk               (video_pll_0_vga_clk_clk),                                            //                   clock.clk
		.reset             (rst_controller_reset_out_reset),                                     //                   reset.reset
		.valid_in          (vga_face_0_avalon_streaming_source_valid),                           //   avalon_streaming_sink.valid
		.startofpacket_in  (vga_face_0_avalon_streaming_source_startofpacket),                   //                        .startofpacket
		.endofpacket_in    (vga_face_0_avalon_streaming_source_endofpacket),                     //                        .endofpacket
		.data_in           (vga_face_0_avalon_streaming_source_data),                            //                        .data
		.ready_out         (vga_face_0_avalon_streaming_source_ready),                           //                        .ready
		.valid_out         (convolution_filter_wrapper_0_avalon_streaming_source_valid),         // avalon_streaming_source.valid
		.startofpacket_out (convolution_filter_wrapper_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.endofpacket_out   (convolution_filter_wrapper_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.data_out          (convolution_filter_wrapper_0_avalon_streaming_source_data),          //                        .data
		.ready_in          (convolution_filter_wrapper_0_avalon_streaming_source_ready),         //                        .ready
		.kernel_select     (kernel_select_kernel_select)                                         //           kernel_select.kernel_select
	);

	pixel_value_filter pixel_value_filter_0 (
		.clk               (video_pll_0_vga_clk_clk),                                            //                   clock.clk
		.reset             (rst_controller_reset_out_reset),                                     //                   reset.reset
		.valid_out         (pixel_value_filter_0_avalon_streaming_source_valid),                 // avalon_streaming_source.valid
		.startofpacket_out (pixel_value_filter_0_avalon_streaming_source_startofpacket),         //                        .startofpacket
		.ready_out         (pixel_value_filter_0_avalon_streaming_source_ready),                 //                        .ready
		.endofpacket_out   (pixel_value_filter_0_avalon_streaming_source_endofpacket),           //                        .endofpacket
		.data_out          (pixel_value_filter_0_avalon_streaming_source_data),                  //                        .data
		.valid_in          (convolution_filter_wrapper_0_avalon_streaming_source_valid),         //   avalon_streaming_sink.valid
		.startofpacket_in  (convolution_filter_wrapper_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.ready_in          (convolution_filter_wrapper_0_avalon_streaming_source_ready),         //                        .ready
		.endofpacket_in    (convolution_filter_wrapper_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.data_in           (convolution_filter_wrapper_0_avalon_streaming_source_data),          //                        .data
		.filter_select     (filter_select_filter_select),                                        //           filter_select.filter_select
		.intensity         (intensity_intensity)                                                 //               intensity.intensity
	);

	vga_face vga_face_0 (
		.clk           (video_pll_0_vga_clk_clk),                          //                   clock.clk
		.reset         (rst_controller_reset_out_reset),                   //                   reset.reset
		.data          (vga_face_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.endofpacket   (vga_face_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.ready         (vga_face_0_avalon_streaming_source_ready),         //                        .ready
		.startofpacket (vga_face_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.valid         (vga_face_0_avalon_streaming_source_valid)          //                        .valid
	);

	vga_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)      // reset_source.reset
	);

	vga_video_vga_controller_0 video_vga_controller_0 (
		.clk           (video_pll_0_vga_clk_clk),                                    //                clk.clk
		.reset         (rst_controller_reset_out_reset),                             //              reset.reset
		.data          (pixel_value_filter_0_avalon_streaming_source_data),          //    avalon_vga_sink.data
		.startofpacket (pixel_value_filter_0_avalon_streaming_source_startofpacket), //                   .startofpacket
		.endofpacket   (pixel_value_filter_0_avalon_streaming_source_endofpacket),   //                   .endofpacket
		.valid         (pixel_value_filter_0_avalon_streaming_source_valid),         //                   .valid
		.ready         (pixel_value_filter_0_avalon_streaming_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                                    // external_interface.export
		.VGA_HS        (vga_HS),                                                     //                   .export
		.VGA_VS        (vga_VS),                                                     //                   .export
		.VGA_BLANK     (vga_BLANK),                                                  //                   .export
		.VGA_SYNC      (vga_SYNC),                                                   //                   .export
		.VGA_R         (vga_R),                                                      //                   .export
		.VGA_G         (vga_G),                                                      //                   .export
		.VGA_B         (vga_B)                                                       //                   .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (video_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
